module saturn_alu (
    i_clk,
    i_reset,
	i_en_alu_prep,
	i_en_alu_calc,
	i_en_alu_save
);

input   wire        i_clk;
input   wire        i_reset;
input   wire    	i_en_alu_prep;
input   wire    	i_en_alu_calc;
input   wire    	i_en_alu_save;


endmodule
