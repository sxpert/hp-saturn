/*
    (c) Raphaël Jacquot 2019
    
		This file is part of hp_saturn.

    hp_saturn is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    any later version.

    hp_saturn is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with Foobar.  If not, see <https://www.gnu.org/licenses/>.

 */

`default_nettype none

`include "saturn_def_alu.v"

module saturn_inst_decoder (
    i_clk,
    i_clk_en,
    i_reset,
    i_phases,
    i_phase,
    i_cycle_ctr,
    
    i_bus_busy,

    i_nibble,
    i_reg_p,
    i_current_pc,

    o_instr_pc,

    o_alu_reg_dest,
    o_alu_reg_src_1,
    o_alu_reg_src_2,
    o_alu_imm_value,
    o_alu_opcode,

    o_jump_length,

    o_instr_type,
    o_instr_decoded,
    o_instr_execute,

    /* debugger interface */
    o_dbg_inst_addr
);

input  wire [0:0]  i_clk;
input  wire [0:0]  i_clk_en;
input  wire [0:0]  i_reset;
input  wire [3:0]  i_phases;
input  wire [1:0]  i_phase;
input  wire [31:0] i_cycle_ctr;

input  wire [0:0]  i_bus_busy;

input  wire [3:0]  i_nibble;
input  wire [3:0]  i_reg_p;
input  wire [19:0] i_current_pc;

output reg  [19:0] o_instr_pc;

output reg  [4:0]  o_alu_reg_dest;
output reg  [4:0]  o_alu_reg_src_1;
output reg  [4:0]  o_alu_reg_src_2;
output reg  [3:0]  o_alu_imm_value;
output reg  [4:0]  o_alu_opcode;

output reg  [2:0]  o_jump_length;

output reg  [3:0]  o_instr_type;
/* instruction is fully decoded */
output reg  [0:0]  o_instr_decoded;
/* instruction is sufficiently decoded to start execution */
output reg  [0:0]  o_instr_execute;

/*
 * debugger interface
 */
/* address of the last instruction */
output reg  [19:0] o_dbg_inst_addr;

/**************************************************************************************************
 *
 * sub-modules go here
 *
 *************************************************************************************************/




/**************************************************************************************************
 *
 * the decoder module
 *
 *************************************************************************************************/

/*
 * process state variables
 */

reg [0:0] just_reset;
reg [0:0] decode_started;

/*
 * decoder block variables
 */

reg [0:0] block_2x;
reg [0:0] block_6x;

/*
 * temporary variables
 */
reg [2:0] jump_counter;

/*
 * initialization
 */

initial begin
    o_alu_reg_dest  = `ALU_REG_NONE;
    o_alu_reg_src_1 = `ALU_REG_NONE;
    o_alu_reg_src_2 = `ALU_REG_NONE;
    o_alu_imm_value = 4'b0;
    o_alu_opcode    = `ALU_OP_NOP;

    o_instr_type    = 4'd15;
    o_instr_decoded = 1'b0;
    o_instr_execute = 1'b0;

    /* debugger interface */
    o_dbg_inst_addr = 20'b0;

    /* internal registers */
    just_reset      = 1'b1;
    decode_started  = 1'b0;

    block_2x        = 1'b0;
    block_6x        = 1'b0;

    /* local variables */
    jump_counter    = 3'd0;
end

/****************************
 *
 * main process
 *
 */

always @(posedge i_clk) begin
  
    /*
     * only do something when nothing is busy doing some other tasks
     * either talking to the bus, or debugging something
     */

    if (i_clk_en && i_bus_busy && i_phases[2] && just_reset) begin
        // $display("DECODER  %0d: [%d] dump registers right after reset", i_phase, i_cycle_ctr);
        just_reset      <= 1'b0;
        o_instr_decoded <= 1'b1;
    end

    if (i_clk_en && !i_bus_busy) begin
 
        if (i_phases[1] && !decode_started) begin
            // $display("DECODER  %0d: [%d] store current PC as instruction start %5h", i_phase, i_cycle_ctr, i_current_pc);
            o_instr_pc   <= i_current_pc;
            /* set the instruction to NOP, to avoid any stray processes */
            o_instr_type <= `INSTR_TYPE_NOP;
        end

        if (i_phases[2] && !decode_started) begin
            $display("DECODER  %0d: [%d] nb= %h - start instruction decoding", i_phase, i_cycle_ctr, i_nibble);

            decode_started <= 1'b1;
            case (i_nibble)
                4'h2: block_2x <= 1'b1;
                4'h6: 
                    begin
                        o_instr_type    <= `INSTR_TYPE_JUMP;
                        o_jump_length   <= 3'd2;
                        jump_counter    <= 3'd0;
                        o_instr_execute <= 1'b1;
                        block_6x        <= 1'b1;
                    end
                default: o_instr_type <= `INSTR_TYPE_NOP;
            endcase
        end

        if (i_phases[2] && decode_started) begin
            $display("DECODER  %0d: [%d] nb= %h - decoding", i_phase, i_cycle_ctr, i_nibble);

            if (block_2x) begin
                $display("DECODER  %0d: [%d] P= %h", i_phase, i_cycle_ctr, i_nibble);
                o_alu_reg_dest  <= `ALU_REG_P;
                o_alu_reg_src_1 <= `ALU_REG_IMM;
                o_alu_reg_src_2 <= `ALU_REG_NONE;
                o_alu_imm_value <= i_nibble;
                o_alu_opcode    <= `ALU_OP_COPY;
                o_instr_type    <= `INSTR_TYPE_ALU;
                o_instr_decoded <= 1'b1;
                o_instr_execute <= 1'b1;
                block_2x        <= 1'b0;
                decode_started  <= 1'b0;
            end

            if (block_6x) begin
                // $display("DECODER  %0d: [%d] GOTO %h", i_phase, i_cycle_ctr, i_nibble);
                jump_counter <= jump_counter + 3'd1;
                if (jump_counter == o_jump_length) begin
                    block_6x        <= 1'b0;
                    o_instr_decoded <= 1'b1;
                    decode_started  <= 1'b0;
                end
            end

        end

        if (i_phases[3]) begin
            // $display("DECODER  %0d: [%d] decoder cleanup", i_phase, i_cycle_ctr);
            o_instr_decoded <= 1'b0;
            o_instr_execute <= 1'b0;
        end

    end


    if (i_reset) begin
        /* stuff that needs reset */
        o_alu_reg_dest  <= `ALU_REG_NONE;
        o_alu_reg_src_1 <= `ALU_REG_NONE;
        o_alu_reg_src_2 <= `ALU_REG_NONE;
        o_alu_imm_value <= 4'b0;
        o_alu_opcode    <= `ALU_OP_NOP;

        o_instr_type    <= 4'd15;
        o_instr_decoded <= 1'b0;
        o_instr_execute <= 1'b0;

        /* debugger interface */
        o_dbg_inst_addr <= 20'b0;

        /* internal registers */
        just_reset      <= 1'b1;
        decode_started  <= 1'b0;

        block_2x        <= 1'b0;
        block_6x        <= 1'b0;

        /* local variables */
        jump_counter    = 3'd0;
    end

end


endmodule
